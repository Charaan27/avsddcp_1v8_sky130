* ========================================= *
* IP Core Name: avsddcp_3V3                 *
* Tech Node: 130nm                          *
* PDK : Sky130 PDK by Google SkyWater	    *
* Name of the author : Charaan S            *
* Company : VLSI System Design Corporation  * 
* ========================================= *


* === INCLUDING SKY130 PDK LIBRARY FILES USING .lib FUNCTION === *
.lib "sky130_fd_pr/models/sky130.lib.spice" tt


* === SKY130 NMOS MODELS === *
xm1 in in v1 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm2 v1 v1 v2 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm3 v2 v2 v3 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm4 v3 v3 v4 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm5 v4 v4 out gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18


* === SKY130 CAPACITOR MODELS === *
xc1  v1 clk1 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xc2  v2 clk2 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xc3  v3 clk1 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xc4  v4 clk2 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xcout1  out gnd sky130_fd_pr__cap_mim_m3_1 w=1 l=100


* === SKY130 RESISTOR MODEL === *
xr1  out gnd gnd sky130_fd_pr__res_high_po_0p69 l=100000


* === CLOCK PULSES (FREQ = 2MHz, Vih = 3.6V(Vih = Vdd+0.3) === *
v2  clk1 gnd pulse(0 3.6 250n 0 0 250n 500n)
v3  clk2 gnd pulse(0 3.6 0 0 0 250n 500n)


* === DC VOLTAGE SOURCE (V=3.3V) === *
v1 in gnd  dc 3.3


* u1  out plot_v1

* === TRANSIENT ANALYSIS STARTS === *
.tran 10e-09 10000e-09 0e-00

.TITLE avsddcp_3V3_cp_out 

* === CONTROL STATEMENTS === * 

.control
run



print allv > plot_data_vclk1.txt
print alli > plot_data_iclk1.txt


* === CHANGING PLOT STYLES === *
set xbrushwidth = 3


* === PLOTTING CLOCKS === *
plot v(clk1) v(clk2)+4


.endc
.end
