magic
tech sky130A
timestamp 1628868665
<< nmos >>
rect 0 2 18 102
rect 154 1 172 101
rect 307 -1 325 99
rect 473 -1 491 99
rect 621 -1 639 99
<< ndiff >>
rect -45 60 0 102
rect -45 42 -32 60
rect -14 42 0 60
rect -45 2 0 42
rect 18 60 63 102
rect 18 42 32 60
rect 50 42 63 60
rect 18 2 63 42
rect 109 59 154 101
rect 109 41 122 59
rect 140 41 154 59
rect 109 1 154 41
rect 172 59 217 101
rect 172 41 186 59
rect 204 41 217 59
rect 172 1 217 41
rect 262 57 307 99
rect 262 39 275 57
rect 293 39 307 57
rect 262 -1 307 39
rect 325 57 370 99
rect 325 39 339 57
rect 357 39 370 57
rect 325 -1 370 39
rect 428 57 473 99
rect 428 39 441 57
rect 459 39 473 57
rect 428 -1 473 39
rect 491 57 536 99
rect 491 39 505 57
rect 523 39 536 57
rect 491 -1 536 39
rect 576 57 621 99
rect 576 39 589 57
rect 607 39 621 57
rect 576 -1 621 39
rect 639 57 684 99
rect 639 39 653 57
rect 671 39 684 57
rect 639 -1 684 39
<< ndiffc >>
rect -32 42 -14 60
rect 32 42 50 60
rect 122 41 140 59
rect 186 41 204 59
rect 275 39 293 57
rect 339 39 357 57
rect 441 39 459 57
rect 505 39 523 57
rect 589 39 607 57
rect 653 39 671 57
<< psubdiff >>
rect 1207 -369 1250 -316
rect 1207 -387 1219 -369
rect 1237 -387 1250 -369
rect 1207 -427 1250 -387
<< psubdiffcont >>
rect 1219 -387 1237 -369
<< poly >>
rect -8 153 26 161
rect -8 135 0 153
rect 18 135 26 153
rect -8 127 26 135
rect 146 152 180 160
rect 146 134 154 152
rect 172 134 180 152
rect 0 102 18 127
rect 146 126 180 134
rect 299 150 333 158
rect 299 132 307 150
rect 325 132 333 150
rect 154 101 172 126
rect 299 124 333 132
rect 465 150 499 158
rect 465 132 473 150
rect 491 132 499 150
rect 465 124 499 132
rect 613 150 647 158
rect 613 132 621 150
rect 639 132 647 150
rect 613 124 647 132
rect 0 -23 18 2
rect 307 99 325 124
rect 473 99 491 124
rect 621 99 639 124
rect 154 -24 172 1
rect 307 -26 325 -1
rect 473 -26 491 -1
rect 621 -26 639 -1
<< polycont >>
rect 0 135 18 153
rect 154 134 172 152
rect 307 132 325 150
rect 473 132 491 150
rect 621 132 639 150
<< locali >>
rect 1267 252 1329 253
rect -98 212 212 233
rect -98 68 -58 212
rect -8 153 58 161
rect 180 160 212 212
rect -8 135 0 153
rect 18 135 58 153
rect -8 127 58 135
rect -98 60 -6 68
rect -98 42 -32 60
rect -14 42 -6 60
rect -98 34 -6 42
rect 24 60 58 127
rect 146 152 212 160
rect 146 134 154 152
rect 172 134 212 152
rect 146 126 212 134
rect 24 42 32 60
rect 50 42 58 60
rect 24 34 58 42
rect 80 59 148 67
rect 80 41 122 59
rect 140 41 148 59
rect -98 -349 -58 34
rect 80 33 148 41
rect 178 59 212 126
rect 178 41 186 59
rect 204 41 212 59
rect 178 33 212 41
rect 231 229 1329 252
rect 231 65 255 229
rect 499 158 531 229
rect 299 150 365 158
rect 299 132 307 150
rect 325 132 365 150
rect 299 124 365 132
rect 465 150 531 158
rect 465 132 473 150
rect 491 132 531 150
rect 465 124 531 132
rect 231 57 301 65
rect 231 39 275 57
rect 293 39 301 57
rect 80 -37 97 33
rect 231 31 301 39
rect 331 57 365 124
rect 331 39 339 57
rect 357 39 365 57
rect 331 31 365 39
rect 392 57 467 65
rect 392 39 441 57
rect 459 39 467 57
rect 392 31 467 39
rect 497 57 531 124
rect 497 39 505 57
rect 523 39 531 57
rect 497 31 531 39
rect 551 192 809 210
rect 551 65 573 192
rect 613 150 679 158
rect 613 132 621 150
rect 639 132 679 150
rect 613 124 679 132
rect 551 57 615 65
rect 551 39 589 57
rect 607 39 615 57
rect 551 31 615 39
rect 645 57 679 124
rect 645 39 653 57
rect 671 39 679 57
rect 331 -37 366 31
rect 80 -54 366 -37
rect 392 -34 424 31
rect 645 -34 679 39
rect 392 -54 679 -34
rect 330 -343 359 -54
rect 645 -115 679 -54
rect 753 -63 809 192
rect 836 -63 884 -15
rect 753 -102 884 -63
rect 520 -145 679 -115
rect 710 -141 1131 -140
rect 1267 -141 1329 229
rect -98 -393 153 -349
rect 330 -387 433 -343
rect 520 -459 564 -145
rect 710 -163 1329 -141
rect 590 -401 638 -334
rect 710 -401 736 -163
rect 1095 -164 1329 -163
rect 590 -435 736 -401
rect 814 -459 862 -336
rect 1211 -369 1245 -361
rect 1211 -387 1219 -369
rect 1237 -387 1245 -369
rect 1211 -395 1245 -387
rect 520 -493 862 -459
<< metal3 >>
rect 819 2 947 130
rect 902 -58 947 2
rect 88 -332 216 -204
rect 368 -326 496 -198
rect 573 -317 701 -189
rect 171 -392 216 -332
rect 451 -386 496 -326
rect 656 -377 701 -317
rect 797 -319 925 -191
rect 880 -379 925 -319
<< mimcap >>
rect 833 61 933 116
rect 833 26 843 61
rect 878 26 933 61
rect 833 16 933 26
rect 102 -273 202 -218
rect 102 -308 112 -273
rect 147 -308 202 -273
rect 102 -318 202 -308
rect 382 -267 482 -212
rect 382 -302 392 -267
rect 427 -302 482 -267
rect 382 -312 482 -302
rect 587 -258 687 -203
rect 587 -293 597 -258
rect 632 -293 687 -258
rect 587 -303 687 -293
rect 811 -260 911 -205
rect 811 -295 821 -260
rect 856 -295 911 -260
rect 811 -305 911 -295
<< mimcapcontact >>
rect 843 26 878 61
rect 112 -308 147 -273
rect 392 -302 427 -267
rect 597 -293 632 -258
rect 821 -295 856 -260
<< metal4 >>
rect 838 61 883 69
rect 838 26 843 61
rect 878 26 883 61
rect 838 -58 883 26
rect 592 -258 637 -250
rect 107 -273 152 -265
rect 107 -308 112 -273
rect 147 -308 152 -273
rect 107 -392 152 -308
rect 387 -267 432 -259
rect 387 -302 392 -267
rect 427 -302 432 -267
rect 387 -386 432 -302
rect 592 -293 597 -258
rect 632 -293 637 -258
rect 592 -377 637 -293
rect 816 -260 861 -252
rect 816 -295 821 -260
rect 856 -295 861 -260
rect 816 -379 861 -295
<< labels >>
rlabel metal4 127 -391 127 -391 5 top
rlabel metal3 192 -391 192 -391 5 bot
rlabel metal4 407 -385 407 -385 5 top
rlabel metal3 472 -385 472 -385 5 bot
rlabel metal3 677 -376 677 -376 5 bot
rlabel metal4 612 -376 612 -376 5 top
rlabel metal3 901 -378 901 -378 5 bot
rlabel metal4 836 -378 836 -378 5 top
rlabel metal3 923 -57 923 -57 5 bot
rlabel metal4 858 -57 858 -57 5 top
<< end >>
